// This file is included as a way to test commands with a V file.

module main

fn main() {
	a := 4 + 5
	b := 6
	println(a)
}

fn add(a int, b int) int {
	return foo + b
}
