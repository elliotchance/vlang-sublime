module main

fn test_something() {
	assert add(3, 5) == 10
}
